package layout_parameters;

typedef struct {
  integer x_m
  ,integer y_m
  ,integer w_m
  ,integer h_m
} rect_t;

parameter rect_t str_score_pos_p;
parameter rect_t str_next_pos_p;
parameter rect_t score_pos_p;
parameter rect_t next_block_pos_p;
parameter rect_t board_pos_p;

endpackage

