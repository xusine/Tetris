module memory_str_score#(
  parameter integer width_p
  ,parameter integer depth_p
)(
  input [$clog2(depth_p)-1:0] addr_i
  ,output logic [width_p-1:0] data_o
);
always_comb unique case(addr_i)
  0: data_o = 0;
  1: data_o = 0;
  2: data_o = 0;
  3: data_o = 0;
  4: data_o = 0;
  5: data_o = 0;
  6: data_o = 0;
  7: data_o = 0;
  8: data_o = 0;
  9: data_o = 0;
  10: data_o = 0;
  11: data_o = 2143289855;
  12: data_o = 2143289855;
  13: data_o = 264241662;
  14: data_o = 264242172;
  15: data_o = 266339324;
  16: data_o = 266339324;
  17: data_o = 266339324;
  18: data_o = 266340348;
  19: data_o = 266340348;
  20: data_o = 267388924;
  21: data_o = 267388924;
  22: data_o = 267390972;
  23: data_o = 267390972;
  24: data_o = 267915260;
  25: data_o = 267915260;
  26: data_o = 267919356;
  27: data_o = 267919356;
  28: data_o = 268181244;
  29: data_o = 268181244;
  30: data_o = 251412220;
  31: data_o = 251412220;
  32: data_o = 251411708;
  33: data_o = 251542780;
  34: data_o = 243154172;
  35: data_o = 243170556;
  36: data_o = 243169532;
  37: data_o = 243235068;
  38: data_o = 239040764;
  39: data_o = 239073532;
  40: data_o = 239071484;
  41: data_o = 239071484;
  42: data_o = 239071484;
  43: data_o = 236974332;
  44: data_o = 236970236;
  45: data_o = 236970236;
  46: data_o = 236970236;
  47: data_o = 235921660;
  48: data_o = 235913468;
  49: data_o = 235913468;
  50: data_o = 235913468;
  51: data_o = 235389180;
  52: data_o = 252150270;
  53: data_o = 2143784959;
  54: data_o = 2143784959;
  55: data_o = 0;
  56: data_o = 0;
  57: data_o = 0;
  58: data_o = 0;
  59: data_o = 0;
  60: data_o = 0;
  61: data_o = 0;
  62: data_o = 0;
  63: data_o = 0;
  64: data_o = 0;
  65: data_o = 0;
  66: data_o = 0;
  67: data_o = 0;
  68: data_o = 0;
  69: data_o = 0;
  70: data_o = 0;
  71: data_o = 0;
  72: data_o = 0;
  73: data_o = 0;
  74: data_o = 0;
  75: data_o = 0;
  76: data_o = 0;
  77: data_o = 0;
  78: data_o = 0;
  79: data_o = 0;
  80: data_o = 0;
  81: data_o = 0;
  82: data_o = 0;
  83: data_o = 0;
  84: data_o = 0;
  85: data_o = 0;
  86: data_o = 0;
  87: data_o = 0;
  88: data_o = 0;
  89: data_o = 536813567;
  90: data_o = 536813567;
  91: data_o = 66585592;
  92: data_o = 33030640;
  93: data_o = 33030624;
  94: data_o = 33031136;
  95: data_o = 16516032;
  96: data_o = 16516032;
  97: data_o = 16517056;
  98: data_o = 8259456;
  99: data_o = 8259456;
  100: data_o = 4067200;
  101: data_o = 4132608;
  102: data_o = 4132608;
  103: data_o = 2039552;
  104: data_o = 2072064;
  105: data_o = 1023488;
  106: data_o = 1048064;
  107: data_o = 1047552;
  108: data_o = 523264;
  109: data_o = 523264;
  110: data_o = 260096;
  111: data_o = 260096;
  112: data_o = 260096;
  113: data_o = 126976;
  114: data_o = 126976;
  115: data_o = 126976;
  116: data_o = 122880;
  117: data_o = 122880;
  118: data_o = 253952;
  119: data_o = 245760;
  120: data_o = 507904;
  121: data_o = 65519616;
  122: data_o = 134184960;
  123: data_o = 134152192;
  124: data_o = 134152192;
  125: data_o = 134086656;
  126: data_o = 66584576;
  127: data_o = 0;
  128: data_o = 0;
  129: data_o = 0;
  130: data_o = 0;
  131: data_o = 0;
  132: data_o = 0;
  133: data_o = 0;
  134: data_o = 0;
  135: data_o = 0;
  136: data_o = 0;
  137: data_o = 0;
  138: data_o = 0;
  139: data_o = 0;
  140: data_o = 0;
  141: data_o = 0;
  142: data_o = 0;
  143: data_o = 0;
  144: data_o = 0;
  145: data_o = 0;
  146: data_o = 0;
  147: data_o = 0;
  148: data_o = 0;
  149: data_o = 0;
  150: data_o = 0;
  151: data_o = 0;
  152: data_o = 0;
  153: data_o = 0;
  154: data_o = 0;
  155: data_o = 0;
  156: data_o = 0;
  157: data_o = 0;
  158: data_o = 0;
  159: data_o = 0;
  160: data_o = 0;
  161: data_o = 0;
  162: data_o = 0;
  163: data_o = 0;
  164: data_o = 0;
  165: data_o = 0;
  166: data_o = 0;
  167: data_o = 0;
  168: data_o = 0;
  169: data_o = 0;
  170: data_o = 0;
  171: data_o = 0;
  172: data_o = 0;
  173: data_o = 0;
  174: data_o = 0;
  175: data_o = 0;
  176: data_o = 0;
  177: data_o = 0;
  178: data_o = 0;
  179: data_o = 0;
  180: data_o = 0;
  181: data_o = 0;
  182: data_o = 0;
  183: data_o = 0;
  184: data_o = 0;
  185: data_o = 0;
  186: data_o = 0;
  187: data_o = 0;
  188: data_o = 0;
  189: data_o = 0;
  190: data_o = 0;
  191: data_o = 0;
  192: data_o = 0;
  193: data_o = 0;
  194: data_o = 0;
  195: data_o = 0;
  196: data_o = 0;
  197: data_o = 0;
  198: data_o = 0;
  199: data_o = 0;
  200: data_o = 0;
  201: data_o = 0;
  202: data_o = 0;
  203: data_o = 1046528;
  204: data_o = 8388464;
  205: data_o = 16777200;
  206: data_o = 33300464;
  207: data_o = 66586608;
  208: data_o = 133170168;
  209: data_o = 132121080;
  210: data_o = 266338552;
  211: data_o = 264241400;
  212: data_o = 264241272;
  213: data_o = 264241272;
  214: data_o = 264241152;
  215: data_o = 264241152;
  216: data_o = 266338304;
  217: data_o = 267386880;
  218: data_o = 133693440;
  219: data_o = 134086656;
  220: data_o = 67076096;
  221: data_o = 33546240;
  222: data_o = 16775168;
  223: data_o = 8388096;
  224: data_o = 2096896;
  225: data_o = 524224;
  226: data_o = 131040;
  227: data_o = 32752;
  228: data_o = 8176;
  229: data_o = 4088;
  230: data_o = 2040;
  231: data_o = 1020;
  232: data_o = 508;
  233: data_o = 503316732;
  234: data_o = 503316732;
  235: data_o = 503316732;
  236: data_o = 520093948;
  237: data_o = 251658492;
  238: data_o = 260047100;
  239: data_o = 260047352;
  240: data_o = 264241656;
  241: data_o = 266339312;
  242: data_o = 267388912;
  243: data_o = 268312544;
  244: data_o = 134217664;
  245: data_o = 127926144;
  246: data_o = 117963776;
  247: data_o = 0;
  248: data_o = 0;
  249: data_o = 0;
  250: data_o = 0;
  251: data_o = 0;
  252: data_o = 0;
  253: data_o = 0;
  254: data_o = 0;
  255: data_o = 0;
  256: data_o = 0;
  257: data_o = 0;
  258: data_o = 0;
  259: data_o = 0;
  260: data_o = 0;
  261: data_o = 0;
  262: data_o = 0;
  263: data_o = 0;
  264: data_o = 0;
  265: data_o = 0;
  266: data_o = 0;
  267: data_o = 0;
  268: data_o = 0;
  269: data_o = 0;
  270: data_o = 0;
  271: data_o = 0;
  272: data_o = 0;
  273: data_o = 0;
  274: data_o = 0;
  275: data_o = 0;
  276: data_o = 0;
  277: data_o = 0;
  278: data_o = 0;
  279: data_o = 0;
  280: data_o = 0;
  281: data_o = 523776;
  282: data_o = 2097024;
  283: data_o = 8388544;
  284: data_o = 16715744;
  285: data_o = 33424368;
  286: data_o = 33293296;
  287: data_o = 66585584;
  288: data_o = 133170160;
  289: data_o = 132121584;
  290: data_o = 132121056;
  291: data_o = 266338304;
  292: data_o = 264241152;
  293: data_o = 264241152;
  294: data_o = 264241152;
  295: data_o = 264241152;
  296: data_o = 264241152;
  297: data_o = 264241152;
  298: data_o = 264241152;
  299: data_o = 264241152;
  300: data_o = 264241152;
  301: data_o = 132120636;
  302: data_o = 132120636;
  303: data_o = 133169276;
  304: data_o = 66060408;
  305: data_o = 66584824;
  306: data_o = 33292784;
  307: data_o = 16713696;
  308: data_o = 8388544;
  309: data_o = 4194176;
  310: data_o = 523776;
  311: data_o = 0;
  312: data_o = 0;
  313: data_o = 0;
  314: data_o = 0;
  315: data_o = 0;
  316: data_o = 0;
  317: data_o = 0;
  318: data_o = 0;
  319: data_o = 0;
  320: data_o = 0;
  321: data_o = 0;
  322: data_o = 0;
  323: data_o = 0;
  324: data_o = 0;
  325: data_o = 0;
  326: data_o = 0;
  327: data_o = 0;
  328: data_o = 0;
  329: data_o = 0;
  330: data_o = 0;
  331: data_o = 0;
  332: data_o = 0;
  333: data_o = 0;
  334: data_o = 0;
  335: data_o = 0;
  336: data_o = 0;
  337: data_o = 0;
  338: data_o = 0;
  339: data_o = 0;
  340: data_o = 0;
  341: data_o = 0;
  342: data_o = 0;
  343: data_o = 0;
  344: data_o = 0;
  345: data_o = 1047552;
  346: data_o = 4194048;
  347: data_o = 8388544;
  348: data_o = 16654304;
  349: data_o = 33294320;
  350: data_o = 66061296;
  351: data_o = 133169656;
  352: data_o = 132121080;
  353: data_o = 264241404;
  354: data_o = 264241404;
  355: data_o = 264241406;
  356: data_o = 528482430;
  357: data_o = 528482430;
  358: data_o = 528482430;
  359: data_o = 528482430;
  360: data_o = 528482430;
  361: data_o = 528482430;
  362: data_o = 528482430;
  363: data_o = 528482430;
  364: data_o = 528482430;
  365: data_o = 264241404;
  366: data_o = 264241404;
  367: data_o = 132121084;
  368: data_o = 132121080;
  369: data_o = 66061296;
  370: data_o = 66586608;
  371: data_o = 33431520;
  372: data_o = 16777152;
  373: data_o = 4194048;
  374: data_o = 1047552;
  375: data_o = 0;
  376: data_o = 0;
  377: data_o = 0;
  378: data_o = 0;
  379: data_o = 0;
  380: data_o = 0;
  381: data_o = 0;
  382: data_o = 0;
  383: data_o = 0;
  384: data_o = 0;
  385: data_o = 0;
  386: data_o = 0;
  387: data_o = 0;
  388: data_o = 0;
  389: data_o = 0;
  390: data_o = 0;
  391: data_o = 0;
  392: data_o = 0;
  393: data_o = 0;
  394: data_o = 0;
  395: data_o = 0;
  396: data_o = 0;
  397: data_o = 0;
  398: data_o = 0;
  399: data_o = 0;
  400: data_o = 0;
  401: data_o = 0;
  402: data_o = 0;
  403: data_o = 0;
  404: data_o = 0;
  405: data_o = 0;
  406: data_o = 0;
  407: data_o = 0;
  408: data_o = 4063232;
  409: data_o = 1073612792;
  410: data_o = 1073618940;
  411: data_o = 16662526;
  412: data_o = 8289918;
  413: data_o = 8322174;
  414: data_o = 8384638;
  415: data_o = 8380542;
  416: data_o = 8372284;
  417: data_o = 8372224;
  418: data_o = 8355840;
  419: data_o = 8323072;
  420: data_o = 8323072;
  421: data_o = 8257536;
  422: data_o = 8257536;
  423: data_o = 8257536;
  424: data_o = 8257536;
  425: data_o = 8257536;
  426: data_o = 8257536;
  427: data_o = 8257536;
  428: data_o = 8257536;
  429: data_o = 8257536;
  430: data_o = 8257536;
  431: data_o = 8257536;
  432: data_o = 8257536;
  433: data_o = 8257536;
  434: data_o = 8257536;
  435: data_o = 8257536;
  436: data_o = 16711680;
  437: data_o = 1073741312;
  438: data_o = 1073741312;
  439: data_o = 0;
  440: data_o = 0;
  441: data_o = 0;
  442: data_o = 0;
  443: data_o = 0;
  444: data_o = 0;
  445: data_o = 0;
  446: data_o = 0;
  447: data_o = 0;
  448: data_o = 0;
  449: data_o = 0;
  450: data_o = 0;
  451: data_o = 0;
  452: data_o = 0;
  453: data_o = 0;
  454: data_o = 0;
  455: data_o = 0;
  456: data_o = 0;
  457: data_o = 0;
  458: data_o = 0;
  459: data_o = 0;
  460: data_o = 0;
  461: data_o = 0;
  462: data_o = 0;
  463: data_o = 0;
  464: data_o = 0;
  465: data_o = 0;
  466: data_o = 0;
  467: data_o = 0;
  468: data_o = 0;
  469: data_o = 0;
  470: data_o = 0;
  471: data_o = 0;
  472: data_o = 0;
  473: data_o = 523264;
  474: data_o = 2096896;
  475: data_o = 8388544;
  476: data_o = 16719840;
  477: data_o = 33294320;
  478: data_o = 33031152;
  479: data_o = 66060792;
  480: data_o = 132121080;
  481: data_o = 132121080;
  482: data_o = 132120828;
  483: data_o = 264241404;
  484: data_o = 264241404;
  485: data_o = 264241404;
  486: data_o = 268435452;
  487: data_o = 268435452;
  488: data_o = 268435452;
  489: data_o = 264241152;
  490: data_o = 264241152;
  491: data_o = 264241152;
  492: data_o = 264241152;
  493: data_o = 132120576;
  494: data_o = 132120696;
  495: data_o = 132120696;
  496: data_o = 66060536;
  497: data_o = 66585072;
  498: data_o = 33293280;
  499: data_o = 16715744;
  500: data_o = 8388544;
  501: data_o = 4194048;
  502: data_o = 523264;
  503: data_o = 0;
  504: data_o = 0;
  505: data_o = 0;
  506: data_o = 0;
  507: data_o = 0;
  508: data_o = 0;
  509: data_o = 0;
  510: data_o = 0;
  511: data_o = 0;
  default: data_o = 'X;
endcase
endmodule
