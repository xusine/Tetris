module memory_str_number#(
  parameter integer width_p
  ,parameter integer depth_p
)(
  input [$clog2(depth_p)-1:0] addr_i
  ,output logic [width_p-1:0] data_o
);
always_comb unique case(addr_i)
  0: data_o = 0;
  1: data_o = 0;
  2: data_o = 0;
  3: data_o = 0;
  4: data_o = 0;
  5: data_o = 0;
  6: data_o = 0;
  7: data_o = 0;
  8: data_o = 0;
  9: data_o = 0;
  10: data_o = 0;
  11: data_o = 522240;
  12: data_o = 2096640;
  13: data_o = 8388480;
  14: data_o = 16719808;
  15: data_o = 16519136;
  16: data_o = 33032160;
  17: data_o = 66585584;
  18: data_o = 66061296;
  19: data_o = 133169656;
  20: data_o = 132121080;
  21: data_o = 132120828;
  22: data_o = 264241404;
  23: data_o = 264241404;
  24: data_o = 264241404;
  25: data_o = 264241404;
  26: data_o = 528482430;
  27: data_o = 528482430;
  28: data_o = 528482430;
  29: data_o = 528482430;
  30: data_o = 528482430;
  31: data_o = 528482430;
  32: data_o = 528482430;
  33: data_o = 528482430;
  34: data_o = 528482430;
  35: data_o = 528482430;
  36: data_o = 528482430;
  37: data_o = 528482430;
  38: data_o = 528482430;
  39: data_o = 528482430;
  40: data_o = 264241404;
  41: data_o = 264241404;
  42: data_o = 264241404;
  43: data_o = 264241404;
  44: data_o = 266338556;
  45: data_o = 132121080;
  46: data_o = 132121080;
  47: data_o = 66061296;
  48: data_o = 66585584;
  49: data_o = 33032160;
  50: data_o = 16519104;
  51: data_o = 16719808;
  52: data_o = 4194176;
  53: data_o = 2096640;
  54: data_o = 522240;
  55: data_o = 0;
  56: data_o = 0;
  57: data_o = 0;
  58: data_o = 0;
  59: data_o = 0;
  60: data_o = 0;
  61: data_o = 0;
  62: data_o = 0;
  63: data_o = 0;
  64: data_o = 0;
  65: data_o = 0;
  66: data_o = 0;
  67: data_o = 0;
  68: data_o = 0;
  69: data_o = 0;
  70: data_o = 0;
  71: data_o = 0;
  72: data_o = 0;
  73: data_o = 0;
  74: data_o = 0;
  75: data_o = 28672;
  76: data_o = 61440;
  77: data_o = 126976;
  78: data_o = 520192;
  79: data_o = 33550336;
  80: data_o = 33550336;
  81: data_o = 520192;
  82: data_o = 258048;
  83: data_o = 258048;
  84: data_o = 258048;
  85: data_o = 258048;
  86: data_o = 258048;
  87: data_o = 258048;
  88: data_o = 258048;
  89: data_o = 258048;
  90: data_o = 258048;
  91: data_o = 258048;
  92: data_o = 258048;
  93: data_o = 258048;
  94: data_o = 258048;
  95: data_o = 258048;
  96: data_o = 258048;
  97: data_o = 258048;
  98: data_o = 258048;
  99: data_o = 258048;
  100: data_o = 258048;
  101: data_o = 258048;
  102: data_o = 258048;
  103: data_o = 258048;
  104: data_o = 258048;
  105: data_o = 258048;
  106: data_o = 258048;
  107: data_o = 258048;
  108: data_o = 258048;
  109: data_o = 258048;
  110: data_o = 258048;
  111: data_o = 258048;
  112: data_o = 258048;
  113: data_o = 258048;
  114: data_o = 258048;
  115: data_o = 522240;
  116: data_o = 1047552;
  117: data_o = 33554400;
  118: data_o = 33554400;
  119: data_o = 0;
  120: data_o = 0;
  121: data_o = 0;
  122: data_o = 0;
  123: data_o = 0;
  124: data_o = 0;
  125: data_o = 0;
  126: data_o = 0;
  127: data_o = 0;
  128: data_o = 0;
  129: data_o = 0;
  130: data_o = 0;
  131: data_o = 0;
  132: data_o = 0;
  133: data_o = 0;
  134: data_o = 0;
  135: data_o = 0;
  136: data_o = 0;
  137: data_o = 0;
  138: data_o = 0;
  139: data_o = 1047552;
  140: data_o = 4194176;
  141: data_o = 16777184;
  142: data_o = 33300464;
  143: data_o = 66062320;
  144: data_o = 132121592;
  145: data_o = 132121080;
  146: data_o = 264241660;
  147: data_o = 264241404;
  148: data_o = 266338556;
  149: data_o = 267387132;
  150: data_o = 267387132;
  151: data_o = 267387132;
  152: data_o = 267387132;
  153: data_o = 132121084;
  154: data_o = 504;
  155: data_o = 504;
  156: data_o = 1016;
  157: data_o = 2032;
  158: data_o = 2016;
  159: data_o = 4064;
  160: data_o = 8128;
  161: data_o = 16256;
  162: data_o = 32512;
  163: data_o = 65024;
  164: data_o = 130048;
  165: data_o = 258048;
  166: data_o = 516096;
  167: data_o = 1032192;
  168: data_o = 2064384;
  169: data_o = 4128768;
  170: data_o = 8257536;
  171: data_o = 16515132;
  172: data_o = 33030204;
  173: data_o = 66060348;
  174: data_o = 65011772;
  175: data_o = 132120700;
  176: data_o = 264241400;
  177: data_o = 528482808;
  178: data_o = 536870904;
  179: data_o = 536870904;
  180: data_o = 536870904;
  181: data_o = 536870904;
  182: data_o = 536870904;
  183: data_o = 0;
  184: data_o = 0;
  185: data_o = 0;
  186: data_o = 0;
  187: data_o = 0;
  188: data_o = 0;
  189: data_o = 0;
  190: data_o = 0;
  191: data_o = 0;
  192: data_o = 0;
  193: data_o = 0;
  194: data_o = 0;
  195: data_o = 0;
  196: data_o = 0;
  197: data_o = 0;
  198: data_o = 0;
  199: data_o = 0;
  200: data_o = 0;
  201: data_o = 0;
  202: data_o = 0;
  203: data_o = 1046528;
  204: data_o = 8388096;
  205: data_o = 16777088;
  206: data_o = 33062848;
  207: data_o = 65019840;
  208: data_o = 62918624;
  209: data_o = 130025440;
  210: data_o = 130025456;
  211: data_o = 132121584;
  212: data_o = 132121584;
  213: data_o = 132121584;
  214: data_o = 132121584;
  215: data_o = 62915568;
  216: data_o = 1008;
  217: data_o = 2016;
  218: data_o = 2016;
  219: data_o = 4032;
  220: data_o = 8128;
  221: data_o = 65280;
  222: data_o = 1048064;
  223: data_o = 1048064;
  224: data_o = 1048320;
  225: data_o = 32704;
  226: data_o = 4064;
  227: data_o = 2032;
  228: data_o = 1008;
  229: data_o = 504;
  230: data_o = 504;
  231: data_o = 252;
  232: data_o = 252;
  233: data_o = 252;
  234: data_o = 65011964;
  235: data_o = 133169404;
  236: data_o = 267387132;
  237: data_o = 267387132;
  238: data_o = 267387388;
  239: data_o = 267387384;
  240: data_o = 266339320;
  241: data_o = 132121584;
  242: data_o = 133171168;
  243: data_o = 66854848;
  244: data_o = 33554304;
  245: data_o = 8388352;
  246: data_o = 2095104;
  247: data_o = 0;
  248: data_o = 0;
  249: data_o = 0;
  250: data_o = 0;
  251: data_o = 0;
  252: data_o = 0;
  253: data_o = 0;
  254: data_o = 0;
  255: data_o = 0;
  256: data_o = 0;
  257: data_o = 0;
  258: data_o = 0;
  259: data_o = 0;
  260: data_o = 0;
  261: data_o = 0;
  262: data_o = 0;
  263: data_o = 0;
  264: data_o = 0;
  265: data_o = 0;
  266: data_o = 0;
  267: data_o = 3968;
  268: data_o = 3968;
  269: data_o = 8064;
  270: data_o = 16256;
  271: data_o = 16256;
  272: data_o = 32640;
  273: data_o = 65408;
  274: data_o = 65408;
  275: data_o = 130944;
  276: data_o = 262016;
  277: data_o = 262016;
  278: data_o = 515968;
  279: data_o = 1023872;
  280: data_o = 1023872;
  281: data_o = 2039680;
  282: data_o = 4071296;
  283: data_o = 4071296;
  284: data_o = 8134528;
  285: data_o = 16260992;
  286: data_o = 16260992;
  287: data_o = 32513920;
  288: data_o = 65019776;
  289: data_o = 65019776;
  290: data_o = 130031488;
  291: data_o = 260054912;
  292: data_o = 260054912;
  293: data_o = 520101760;
  294: data_o = 1040195456;
  295: data_o = 1073741823;
  296: data_o = 1073741823;
  297: data_o = 1073741823;
  298: data_o = 8064;
  299: data_o = 8064;
  300: data_o = 8064;
  301: data_o = 8064;
  302: data_o = 8064;
  303: data_o = 8064;
  304: data_o = 8064;
  305: data_o = 8064;
  306: data_o = 8064;
  307: data_o = 8064;
  308: data_o = 16320;
  309: data_o = 524286;
  310: data_o = 524286;
  311: data_o = 0;
  312: data_o = 0;
  313: data_o = 0;
  314: data_o = 0;
  315: data_o = 0;
  316: data_o = 0;
  317: data_o = 0;
  318: data_o = 0;
  319: data_o = 0;
  320: data_o = 0;
  321: data_o = 0;
  322: data_o = 0;
  323: data_o = 0;
  324: data_o = 0;
  325: data_o = 0;
  326: data_o = 0;
  327: data_o = 0;
  328: data_o = 0;
  329: data_o = 0;
  330: data_o = 0;
  331: data_o = 33554424;
  332: data_o = 33554424;
  333: data_o = 33554424;
  334: data_o = 33554424;
  335: data_o = 33554416;
  336: data_o = 31457280;
  337: data_o = 31457280;
  338: data_o = 31457280;
  339: data_o = 31457280;
  340: data_o = 31457280;
  341: data_o = 31457280;
  342: data_o = 31457280;
  343: data_o = 29360128;
  344: data_o = 62914560;
  345: data_o = 62914560;
  346: data_o = 63438336;
  347: data_o = 65011584;
  348: data_o = 67108800;
  349: data_o = 66985952;
  350: data_o = 66586608;
  351: data_o = 66061296;
  352: data_o = 65012728;
  353: data_o = 65012216;
  354: data_o = 58720760;
  355: data_o = 508;
  356: data_o = 252;
  357: data_o = 252;
  358: data_o = 252;
  359: data_o = 252;
  360: data_o = 252;
  361: data_o = 65011964;
  362: data_o = 133169404;
  363: data_o = 267387132;
  364: data_o = 267387132;
  365: data_o = 267387384;
  366: data_o = 267387384;
  367: data_o = 266338808;
  368: data_o = 266339312;
  369: data_o = 132122608;
  370: data_o = 66064352;
  371: data_o = 33300416;
  372: data_o = 16777088;
  373: data_o = 8388352;
  374: data_o = 1047552;
  375: data_o = 0;
  376: data_o = 0;
  377: data_o = 0;
  378: data_o = 0;
  379: data_o = 0;
  380: data_o = 0;
  381: data_o = 0;
  382: data_o = 0;
  383: data_o = 0;
  384: data_o = 0;
  385: data_o = 0;
  386: data_o = 0;
  387: data_o = 0;
  388: data_o = 0;
  389: data_o = 0;
  390: data_o = 0;
  391: data_o = 0;
  392: data_o = 0;
  393: data_o = 0;
  394: data_o = 0;
  395: data_o = 130816;
  396: data_o = 1048512;
  397: data_o = 2097136;
  398: data_o = 4163568;
  399: data_o = 8258552;
  400: data_o = 16516088;
  401: data_o = 33031160;
  402: data_o = 66061304;
  403: data_o = 65012208;
  404: data_o = 132120576;
  405: data_o = 130023424;
  406: data_o = 130023424;
  407: data_o = 264241152;
  408: data_o = 264241152;
  409: data_o = 264241152;
  410: data_o = 260046848;
  411: data_o = 528743936;
  412: data_o = 530579392;
  413: data_o = 532676576;
  414: data_o = 536809456;
  415: data_o = 536609784;
  416: data_o = 536347128;
  417: data_o = 535822844;
  418: data_o = 534774012;
  419: data_o = 532676860;
  420: data_o = 532676734;
  421: data_o = 528482430;
  422: data_o = 528482430;
  423: data_o = 528482430;
  424: data_o = 528482430;
  425: data_o = 528482430;
  426: data_o = 264241278;
  427: data_o = 264241278;
  428: data_o = 264241278;
  429: data_o = 264241406;
  430: data_o = 132120828;
  431: data_o = 133169404;
  432: data_o = 66060792;
  433: data_o = 66585080;
  434: data_o = 33293296;
  435: data_o = 16715744;
  436: data_o = 8388544;
  437: data_o = 4194176;
  438: data_o = 523264;
  439: data_o = 0;
  440: data_o = 0;
  441: data_o = 0;
  442: data_o = 0;
  443: data_o = 0;
  444: data_o = 0;
  445: data_o = 0;
  446: data_o = 0;
  447: data_o = 0;
  448: data_o = 0;
  449: data_o = 0;
  450: data_o = 0;
  451: data_o = 0;
  452: data_o = 0;
  453: data_o = 0;
  454: data_o = 0;
  455: data_o = 0;
  456: data_o = 0;
  457: data_o = 0;
  458: data_o = 0;
  459: data_o = 67108860;
  460: data_o = 134217724;
  461: data_o = 134217724;
  462: data_o = 134217724;
  463: data_o = 134217720;
  464: data_o = 133169392;
  465: data_o = 130023920;
  466: data_o = 125829600;
  467: data_o = 260047840;
  468: data_o = 251659200;
  469: data_o = 251660224;
  470: data_o = 251662208;
  471: data_o = 3968;
  472: data_o = 7936;
  473: data_o = 7936;
  474: data_o = 15872;
  475: data_o = 15872;
  476: data_o = 32256;
  477: data_o = 31744;
  478: data_o = 64512;
  479: data_o = 63488;
  480: data_o = 129024;
  481: data_o = 129024;
  482: data_o = 126976;
  483: data_o = 258048;
  484: data_o = 258048;
  485: data_o = 520192;
  486: data_o = 516096;
  487: data_o = 516096;
  488: data_o = 516096;
  489: data_o = 1040384;
  490: data_o = 1040384;
  491: data_o = 1040384;
  492: data_o = 1040384;
  493: data_o = 2088960;
  494: data_o = 2088960;
  495: data_o = 2088960;
  496: data_o = 2088960;
  497: data_o = 2088960;
  498: data_o = 2088960;
  499: data_o = 2088960;
  500: data_o = 2088960;
  501: data_o = 2088960;
  502: data_o = 1032192;
  503: data_o = 0;
  504: data_o = 0;
  505: data_o = 0;
  506: data_o = 0;
  507: data_o = 0;
  508: data_o = 0;
  509: data_o = 0;
  510: data_o = 0;
  511: data_o = 0;
  512: data_o = 0;
  513: data_o = 0;
  514: data_o = 0;
  515: data_o = 0;
  516: data_o = 0;
  517: data_o = 0;
  518: data_o = 0;
  519: data_o = 0;
  520: data_o = 0;
  521: data_o = 0;
  522: data_o = 0;
  523: data_o = 1047552;
  524: data_o = 8388480;
  525: data_o = 16777152;
  526: data_o = 33431520;
  527: data_o = 66586608;
  528: data_o = 133170168;
  529: data_o = 132121080;
  530: data_o = 266338812;
  531: data_o = 264241404;
  532: data_o = 264241404;
  533: data_o = 264241404;
  534: data_o = 264241404;
  535: data_o = 266338556;
  536: data_o = 267387132;
  537: data_o = 133169656;
  538: data_o = 133956088;
  539: data_o = 66978800;
  540: data_o = 67078112;
  541: data_o = 33550272;
  542: data_o = 16777088;
  543: data_o = 4193792;
  544: data_o = 8388352;
  545: data_o = 16777088;
  546: data_o = 33095616;
  547: data_o = 66093024;
  548: data_o = 132128752;
  549: data_o = 266342392;
  550: data_o = 264243192;
  551: data_o = 264242168;
  552: data_o = 532677116;
  553: data_o = 528482812;
  554: data_o = 528482556;
  555: data_o = 528482556;
  556: data_o = 528482556;
  557: data_o = 528482556;
  558: data_o = 532676860;
  559: data_o = 264241656;
  560: data_o = 266338808;
  561: data_o = 132121584;
  562: data_o = 133695472;
  563: data_o = 66854880;
  564: data_o = 16777152;
  565: data_o = 8388352;
  566: data_o = 1047552;
  567: data_o = 0;
  568: data_o = 0;
  569: data_o = 0;
  570: data_o = 0;
  571: data_o = 0;
  572: data_o = 0;
  573: data_o = 0;
  574: data_o = 0;
  575: data_o = 0;
  576: data_o = 0;
  577: data_o = 0;
  578: data_o = 0;
  579: data_o = 0;
  580: data_o = 0;
  581: data_o = 0;
  582: data_o = 0;
  583: data_o = 0;
  584: data_o = 0;
  585: data_o = 0;
  586: data_o = 0;
  587: data_o = 1046528;
  588: data_o = 8388352;
  589: data_o = 16777088;
  590: data_o = 33431488;
  591: data_o = 66586592;
  592: data_o = 133170160;
  593: data_o = 132121072;
  594: data_o = 264241656;
  595: data_o = 264241400;
  596: data_o = 264241404;
  597: data_o = 528482556;
  598: data_o = 528482428;
  599: data_o = 528482428;
  600: data_o = 528482430;
  601: data_o = 528482430;
  602: data_o = 528482430;
  603: data_o = 528482430;
  604: data_o = 528482430;
  605: data_o = 532676862;
  606: data_o = 532676862;
  607: data_o = 264241662;
  608: data_o = 266339326;
  609: data_o = 267388926;
  610: data_o = 133697534;
  611: data_o = 66863102;
  612: data_o = 33554302;
  613: data_o = 16776446;
  614: data_o = 2093308;
  615: data_o = 252;
  616: data_o = 252;
  617: data_o = 252;
  618: data_o = 504;
  619: data_o = 504;
  620: data_o = 504;
  621: data_o = 1008;
  622: data_o = 65012720;
  623: data_o = 133171168;
  624: data_o = 133173216;
  625: data_o = 133173184;
  626: data_o = 133185408;
  627: data_o = 133758720;
  628: data_o = 67108352;
  629: data_o = 33552384;
  630: data_o = 4186112;
  631: data_o = 0;
  632: data_o = 0;
  633: data_o = 0;
  634: data_o = 0;
  635: data_o = 0;
  636: data_o = 0;
  637: data_o = 0;
  638: data_o = 0;
  639: data_o = 0;
  default: data_o = 'X;
endcase
endmodule
