module game_top_logic #(
  parameter integer width_p = 16
  ,parameter integer height_p = 32
)(
  input clk_i
  ,input reset_i

  ,input down_clk_i

  ,input left_i
  ,input right_i
  ,input rotate_i

);


endmodule