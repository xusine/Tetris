module memory_character#(
  parameter integer width_p
  ,parameter integer depth_p
)(
  input [$clog2(depth_p)-1:0] addr_i
  ,output logic [width_p-1:0] data_o
);
always_comb unique case(addr_i)
  0: data_o = 0;
  1: data_o = 0;
  2: data_o = 0;
  3: data_o = 0;
  4: data_o = 0;
  5: data_o = 0;
  6: data_o = 1046528;
  7: data_o = 4193792;
  8: data_o = 8388352;
  9: data_o = 33554304;
  10: data_o = 33554368;
  11: data_o = 66592736;
  12: data_o = 133173216;
  13: data_o = 132122592;
  14: data_o = 264242160;
  15: data_o = 264242160;
  16: data_o = 264242160;
  17: data_o = 264242160;
  18: data_o = 264242160;
  19: data_o = 264241152;
  20: data_o = 264241152;
  21: data_o = 266338304;
  22: data_o = 132120576;
  23: data_o = 133169152;
  24: data_o = 66846720;
  25: data_o = 66977792;
  26: data_o = 33488896;
  27: data_o = 8355840;
  28: data_o = 4186112;
  29: data_o = 2093056;
  30: data_o = 1047552;
  31: data_o = 261888;
  32: data_o = 130944;
  33: data_o = 32704;
  34: data_o = 16352;
  35: data_o = 4080;
  36: data_o = 2032;
  37: data_o = 1016;
  38: data_o = 504;
  39: data_o = 1056965112;
  40: data_o = 1056965112;
  41: data_o = 1056965112;
  42: data_o = 520094200;
  43: data_o = 520094200;
  44: data_o = 528482808;
  45: data_o = 528482808;
  46: data_o = 528483312;
  47: data_o = 264243184;
  48: data_o = 267390944;
  49: data_o = 134217696;
  50: data_o = 67108800;
  51: data_o = 33554304;
  52: data_o = 16776960;
  53: data_o = 4193280;
  54: data_o = 516096;
  55: data_o = 0;
  56: data_o = 0;
  57: data_o = 0;
  58: data_o = 0;
  59: data_o = 0;
  60: data_o = 0;
  61: data_o = 0;
  62: data_o = 0;
  63: data_o = 0;
  64: data_o = 0;
  65: data_o = 0;
  66: data_o = 0;
  67: data_o = 0;
  68: data_o = 0;
  69: data_o = 0;
  70: data_o = 523264;
  71: data_o = 2096896;
  72: data_o = 4194176;
  73: data_o = 8388544;
  74: data_o = 16777152;
  75: data_o = 33294304;
  76: data_o = 33031152;
  77: data_o = 66061296;
  78: data_o = 66060792;
  79: data_o = 132121080;
  80: data_o = 130023928;
  81: data_o = 264241400;
  82: data_o = 264241404;
  83: data_o = 260047100;
  84: data_o = 260047100;
  85: data_o = 528482556;
  86: data_o = 528482556;
  87: data_o = 528482304;
  88: data_o = 528482304;
  89: data_o = 520093696;
  90: data_o = 520093696;
  91: data_o = 520093696;
  92: data_o = 520093696;
  93: data_o = 520093696;
  94: data_o = 520093696;
  95: data_o = 1056964608;
  96: data_o = 520093696;
  97: data_o = 520093696;
  98: data_o = 520093696;
  99: data_o = 520093696;
  100: data_o = 528482556;
  101: data_o = 528482556;
  102: data_o = 528482556;
  103: data_o = 528482556;
  104: data_o = 528482552;
  105: data_o = 260047096;
  106: data_o = 264241656;
  107: data_o = 264241656;
  108: data_o = 132121080;
  109: data_o = 132121584;
  110: data_o = 66061296;
  111: data_o = 66586608;
  112: data_o = 33296352;
  113: data_o = 33554368;
  114: data_o = 16777152;
  115: data_o = 8388480;
  116: data_o = 4194048;
  117: data_o = 1047552;
  118: data_o = 122880;
  119: data_o = 0;
  120: data_o = 0;
  121: data_o = 0;
  122: data_o = 0;
  123: data_o = 0;
  124: data_o = 0;
  125: data_o = 0;
  126: data_o = 0;
  127: data_o = 0;
  128: data_o = 0;
  129: data_o = 0;
  130: data_o = 0;
  131: data_o = 0;
  132: data_o = 0;
  133: data_o = 0;
  134: data_o = 2093056;
  135: data_o = 8387584;
  136: data_o = 16776960;
  137: data_o = 33554304;
  138: data_o = 67108800;
  139: data_o = 66592704;
  140: data_o = 132124640;
  141: data_o = 130025440;
  142: data_o = 264242160;
  143: data_o = 260047856;
  144: data_o = 260047344;
  145: data_o = 528482808;
  146: data_o = 528482808;
  147: data_o = 520094200;
  148: data_o = 520094200;
  149: data_o = 520093944;
  150: data_o = 1056964856;
  151: data_o = 1056964856;
  152: data_o = 1056964860;
  153: data_o = 1056964860;
  154: data_o = 1056964860;
  155: data_o = 1056964860;
  156: data_o = 1056964860;
  157: data_o = 1056964860;
  158: data_o = 1056964860;
  159: data_o = 1056964860;
  160: data_o = 1056964860;
  161: data_o = 1056964860;
  162: data_o = 1056964860;
  163: data_o = 1056964860;
  164: data_o = 1056964856;
  165: data_o = 1056964856;
  166: data_o = 1056964856;
  167: data_o = 520094200;
  168: data_o = 520094200;
  169: data_o = 528482808;
  170: data_o = 528482808;
  171: data_o = 528482800;
  172: data_o = 260047856;
  173: data_o = 264242160;
  174: data_o = 264242144;
  175: data_o = 132122592;
  176: data_o = 133173184;
  177: data_o = 66863040;
  178: data_o = 33554304;
  179: data_o = 16776960;
  180: data_o = 8388096;
  181: data_o = 4192256;
  182: data_o = 507904;
  183: data_o = 0;
  184: data_o = 0;
  185: data_o = 0;
  186: data_o = 0;
  187: data_o = 0;
  188: data_o = 0;
  189: data_o = 0;
  190: data_o = 0;
  191: data_o = 0;
  192: data_o = 0;
  193: data_o = 0;
  194: data_o = 0;
  195: data_o = 0;
  196: data_o = 0;
  197: data_o = 0;
  198: data_o = 536866816;
  199: data_o = 536870400;
  200: data_o = 536870656;
  201: data_o = 536870784;
  202: data_o = 536870848;
  203: data_o = 528490464;
  204: data_o = 528486384;
  205: data_o = 528484336;
  206: data_o = 528483312;
  207: data_o = 528482808;
  208: data_o = 528482808;
  209: data_o = 528482808;
  210: data_o = 528482808;
  211: data_o = 528482808;
  212: data_o = 528482808;
  213: data_o = 528482808;
  214: data_o = 528482808;
  215: data_o = 528483312;
  216: data_o = 528483312;
  217: data_o = 528484336;
  218: data_o = 528490464;
  219: data_o = 536870848;
  220: data_o = 536870784;
  221: data_o = 536870656;
  222: data_o = 536870400;
  223: data_o = 536868864;
  224: data_o = 528546816;
  225: data_o = 528546816;
  226: data_o = 528514048;
  227: data_o = 528514560;
  228: data_o = 528514560;
  229: data_o = 528498432;
  230: data_o = 528498432;
  231: data_o = 528498432;
  232: data_o = 528490368;
  233: data_o = 528490368;
  234: data_o = 528486336;
  235: data_o = 528486336;
  236: data_o = 528486336;
  237: data_o = 528484320;
  238: data_o = 528484320;
  239: data_o = 528483296;
  240: data_o = 528483312;
  241: data_o = 528483312;
  242: data_o = 528482808;
  243: data_o = 528482808;
  244: data_o = 528482808;
  245: data_o = 528482556;
  246: data_o = 528482556;
  247: data_o = 0;
  248: data_o = 0;
  249: data_o = 0;
  250: data_o = 0;
  251: data_o = 0;
  252: data_o = 0;
  253: data_o = 0;
  254: data_o = 0;
  255: data_o = 0;
  256: data_o = 0;
  257: data_o = 0;
  258: data_o = 0;
  259: data_o = 0;
  260: data_o = 0;
  261: data_o = 0;
  262: data_o = 268435440;
  263: data_o = 268435440;
  264: data_o = 268435440;
  265: data_o = 268435440;
  266: data_o = 268435440;
  267: data_o = 264241152;
  268: data_o = 264241152;
  269: data_o = 264241152;
  270: data_o = 264241152;
  271: data_o = 264241152;
  272: data_o = 264241152;
  273: data_o = 264241152;
  274: data_o = 264241152;
  275: data_o = 264241152;
  276: data_o = 264241152;
  277: data_o = 264241152;
  278: data_o = 264241152;
  279: data_o = 264241152;
  280: data_o = 264241152;
  281: data_o = 264241152;
  282: data_o = 268435424;
  283: data_o = 268435424;
  284: data_o = 268435424;
  285: data_o = 268435424;
  286: data_o = 268435424;
  287: data_o = 264241152;
  288: data_o = 264241152;
  289: data_o = 264241152;
  290: data_o = 264241152;
  291: data_o = 264241152;
  292: data_o = 264241152;
  293: data_o = 264241152;
  294: data_o = 264241152;
  295: data_o = 264241152;
  296: data_o = 264241152;
  297: data_o = 264241152;
  298: data_o = 264241152;
  299: data_o = 264241152;
  300: data_o = 264241152;
  301: data_o = 264241152;
  302: data_o = 264241152;
  303: data_o = 264241152;
  304: data_o = 264241152;
  305: data_o = 264241152;
  306: data_o = 268435448;
  307: data_o = 268435448;
  308: data_o = 268435448;
  309: data_o = 268435448;
  310: data_o = 268435448;
  311: data_o = 0;
  312: data_o = 0;
  313: data_o = 0;
  314: data_o = 0;
  315: data_o = 0;
  316: data_o = 0;
  317: data_o = 0;
  318: data_o = 0;
  319: data_o = 0;
  320: data_o = 0;
  321: data_o = 0;
  322: data_o = 0;
  323: data_o = 0;
  324: data_o = 0;
  325: data_o = 0;
  326: data_o = 532677112;
  327: data_o = 532677112;
  328: data_o = 534774264;
  329: data_o = 534774264;
  330: data_o = 534774264;
  331: data_o = 535822840;
  332: data_o = 535822840;
  333: data_o = 536347128;
  334: data_o = 536347128;
  335: data_o = 536347128;
  336: data_o = 536609272;
  337: data_o = 536609272;
  338: data_o = 536609272;
  339: data_o = 536740344;
  340: data_o = 532546040;
  341: data_o = 532546040;
  342: data_o = 532611576;
  343: data_o = 530514424;
  344: data_o = 530514424;
  345: data_o = 530547192;
  346: data_o = 529498616;
  347: data_o = 529498616;
  348: data_o = 529515000;
  349: data_o = 528990712;
  350: data_o = 528998904;
  351: data_o = 528736760;
  352: data_o = 528736760;
  353: data_o = 528740856;
  354: data_o = 528609784;
  355: data_o = 528609784;
  356: data_o = 528611832;
  357: data_o = 528546296;
  358: data_o = 528546296;
  359: data_o = 528547320;
  360: data_o = 528514552;
  361: data_o = 528514552;
  362: data_o = 528515064;
  363: data_o = 528498680;
  364: data_o = 528498680;
  365: data_o = 528498680;
  366: data_o = 528490488;
  367: data_o = 528490488;
  368: data_o = 528486392;
  369: data_o = 528486392;
  370: data_o = 528486392;
  371: data_o = 528484344;
  372: data_o = 528484344;
  373: data_o = 528484344;
  374: data_o = 528483320;
  375: data_o = 0;
  376: data_o = 0;
  377: data_o = 0;
  378: data_o = 0;
  379: data_o = 0;
  380: data_o = 0;
  381: data_o = 0;
  382: data_o = 0;
  383: data_o = 0;
  384: data_o = 0;
  385: data_o = 0;
  386: data_o = 0;
  387: data_o = 0;
  388: data_o = 0;
  389: data_o = 0;
  390: data_o = 268435440;
  391: data_o = 268435440;
  392: data_o = 268435440;
  393: data_o = 268435440;
  394: data_o = 268435440;
  395: data_o = 264241152;
  396: data_o = 264241152;
  397: data_o = 264241152;
  398: data_o = 264241152;
  399: data_o = 264241152;
  400: data_o = 264241152;
  401: data_o = 264241152;
  402: data_o = 264241152;
  403: data_o = 264241152;
  404: data_o = 264241152;
  405: data_o = 264241152;
  406: data_o = 264241152;
  407: data_o = 264241152;
  408: data_o = 264241152;
  409: data_o = 264241152;
  410: data_o = 268435424;
  411: data_o = 268435424;
  412: data_o = 268435424;
  413: data_o = 268435424;
  414: data_o = 268435424;
  415: data_o = 264241152;
  416: data_o = 264241152;
  417: data_o = 264241152;
  418: data_o = 264241152;
  419: data_o = 264241152;
  420: data_o = 264241152;
  421: data_o = 264241152;
  422: data_o = 264241152;
  423: data_o = 264241152;
  424: data_o = 264241152;
  425: data_o = 264241152;
  426: data_o = 264241152;
  427: data_o = 264241152;
  428: data_o = 264241152;
  429: data_o = 264241152;
  430: data_o = 264241152;
  431: data_o = 264241152;
  432: data_o = 264241152;
  433: data_o = 264241152;
  434: data_o = 268435448;
  435: data_o = 268435448;
  436: data_o = 268435448;
  437: data_o = 268435448;
  438: data_o = 268435448;
  439: data_o = 0;
  440: data_o = 0;
  441: data_o = 0;
  442: data_o = 0;
  443: data_o = 0;
  444: data_o = 0;
  445: data_o = 0;
  446: data_o = 0;
  447: data_o = 0;
  448: data_o = 0;
  449: data_o = 0;
  450: data_o = 0;
  451: data_o = 0;
  452: data_o = 0;
  453: data_o = 0;
  454: data_o = 528482808;
  455: data_o = 528482800;
  456: data_o = 260047856;
  457: data_o = 264242144;
  458: data_o = 130025440;
  459: data_o = 132122592;
  460: data_o = 132124608;
  461: data_o = 65015744;
  462: data_o = 66064256;
  463: data_o = 32513920;
  464: data_o = 33038080;
  465: data_o = 16269056;
  466: data_o = 16531200;
  467: data_o = 16530944;
  468: data_o = 8158720;
  469: data_o = 8289280;
  470: data_o = 4127744;
  471: data_o = 4192256;
  472: data_o = 2095104;
  473: data_o = 2095104;
  474: data_o = 2093056;
  475: data_o = 1044480;
  476: data_o = 1040384;
  477: data_o = 1040384;
  478: data_o = 1044480;
  479: data_o = 2093056;
  480: data_o = 2095104;
  481: data_o = 2095104;
  482: data_o = 4192256;
  483: data_o = 4127744;
  484: data_o = 8289280;
  485: data_o = 8158720;
  486: data_o = 16547328;
  487: data_o = 16531200;
  488: data_o = 33046272;
  489: data_o = 33038080;
  490: data_o = 32513920;
  491: data_o = 66064256;
  492: data_o = 65015744;
  493: data_o = 132122560;
  494: data_o = 132122592;
  495: data_o = 264243168;
  496: data_o = 264242160;
  497: data_o = 260047856;
  498: data_o = 528482800;
  499: data_o = 520094200;
  500: data_o = 1056964856;
  501: data_o = 1056964860;
  502: data_o = 2113929468;
  503: data_o = 0;
  504: data_o = 0;
  505: data_o = 0;
  506: data_o = 0;
  507: data_o = 0;
  508: data_o = 0;
  509: data_o = 0;
  510: data_o = 0;
  511: data_o = 0;
  512: data_o = 0;
  513: data_o = 0;
  514: data_o = 0;
  515: data_o = 0;
  516: data_o = 0;
  517: data_o = 0;
  518: data_o = 536870904;
  519: data_o = 536870904;
  520: data_o = 536870904;
  521: data_o = 536870904;
  522: data_o = 536870904;
  523: data_o = 516096;
  524: data_o = 516096;
  525: data_o = 516096;
  526: data_o = 516096;
  527: data_o = 516096;
  528: data_o = 516096;
  529: data_o = 516096;
  530: data_o = 516096;
  531: data_o = 516096;
  532: data_o = 516096;
  533: data_o = 516096;
  534: data_o = 516096;
  535: data_o = 516096;
  536: data_o = 516096;
  537: data_o = 516096;
  538: data_o = 516096;
  539: data_o = 516096;
  540: data_o = 516096;
  541: data_o = 516096;
  542: data_o = 516096;
  543: data_o = 516096;
  544: data_o = 516096;
  545: data_o = 516096;
  546: data_o = 516096;
  547: data_o = 516096;
  548: data_o = 516096;
  549: data_o = 516096;
  550: data_o = 516096;
  551: data_o = 516096;
  552: data_o = 516096;
  553: data_o = 516096;
  554: data_o = 516096;
  555: data_o = 516096;
  556: data_o = 516096;
  557: data_o = 516096;
  558: data_o = 516096;
  559: data_o = 516096;
  560: data_o = 516096;
  561: data_o = 516096;
  562: data_o = 516096;
  563: data_o = 516096;
  564: data_o = 516096;
  565: data_o = 516096;
  566: data_o = 516096;
  567: data_o = 0;
  568: data_o = 0;
  569: data_o = 0;
  570: data_o = 0;
  571: data_o = 0;
  572: data_o = 0;
  573: data_o = 0;
  574: data_o = 0;
  575: data_o = 0;
  576: data_o = 0;
  577: data_o = 0;
  578: data_o = 0;
  579: data_o = 0;
  580: data_o = 0;
  581: data_o = 0;
  582: data_o = 1044480;
  583: data_o = 4192256;
  584: data_o = 8388096;
  585: data_o = 16776960;
  586: data_o = 33554304;
  587: data_o = 66600832;
  588: data_o = 66068416;
  589: data_o = 132124608;
  590: data_o = 132122592;
  591: data_o = 264243168;
  592: data_o = 264242160;
  593: data_o = 528483312;
  594: data_o = 528483312;
  595: data_o = 528482808;
  596: data_o = 528482808;
  597: data_o = 520094200;
  598: data_o = 1056965112;
  599: data_o = 1056965112;
  600: data_o = 1056964856;
  601: data_o = 1056964856;
  602: data_o = 1056964856;
  603: data_o = 1056964856;
  604: data_o = 1056964856;
  605: data_o = 1056964856;
  606: data_o = 1056964856;
  607: data_o = 1056964856;
  608: data_o = 1056964856;
  609: data_o = 1056964856;
  610: data_o = 1056964856;
  611: data_o = 1056964856;
  612: data_o = 1056965112;
  613: data_o = 1056965112;
  614: data_o = 520094200;
  615: data_o = 528482808;
  616: data_o = 528482808;
  617: data_o = 528482800;
  618: data_o = 528483312;
  619: data_o = 264242160;
  620: data_o = 264243168;
  621: data_o = 266340320;
  622: data_o = 132124640;
  623: data_o = 133173184;
  624: data_o = 66592640;
  625: data_o = 33324928;
  626: data_o = 16776960;
  627: data_o = 16776704;
  628: data_o = 4193280;
  629: data_o = 2093056;
  630: data_o = 245760;
  631: data_o = 0;
  632: data_o = 0;
  633: data_o = 0;
  634: data_o = 0;
  635: data_o = 0;
  636: data_o = 0;
  637: data_o = 0;
  638: data_o = 0;
  639: data_o = 0;
  640: data_o = 0;
  641: data_o = 0;
  642: data_o = 0;
  643: data_o = 0;
  644: data_o = 0;
  645: data_o = 0;
  646: data_o = 61440;
  647: data_o = 61440;
  648: data_o = 126976;
  649: data_o = 126976;
  650: data_o = 258048;
  651: data_o = 1044480;
  652: data_o = 8384512;
  653: data_o = 67104768;
  654: data_o = 67104768;
  655: data_o = 67104768;
  656: data_o = 258048;
  657: data_o = 258048;
  658: data_o = 258048;
  659: data_o = 258048;
  660: data_o = 258048;
  661: data_o = 258048;
  662: data_o = 258048;
  663: data_o = 258048;
  664: data_o = 258048;
  665: data_o = 258048;
  666: data_o = 258048;
  667: data_o = 258048;
  668: data_o = 258048;
  669: data_o = 258048;
  670: data_o = 258048;
  671: data_o = 258048;
  672: data_o = 258048;
  673: data_o = 258048;
  674: data_o = 258048;
  675: data_o = 258048;
  676: data_o = 258048;
  677: data_o = 258048;
  678: data_o = 258048;
  679: data_o = 258048;
  680: data_o = 258048;
  681: data_o = 258048;
  682: data_o = 258048;
  683: data_o = 258048;
  684: data_o = 258048;
  685: data_o = 258048;
  686: data_o = 258048;
  687: data_o = 258048;
  688: data_o = 258048;
  689: data_o = 258048;
  690: data_o = 258048;
  691: data_o = 258048;
  692: data_o = 258048;
  693: data_o = 258048;
  694: data_o = 258048;
  695: data_o = 0;
  696: data_o = 0;
  697: data_o = 0;
  698: data_o = 0;
  699: data_o = 0;
  700: data_o = 0;
  701: data_o = 0;
  702: data_o = 0;
  703: data_o = 0;
  704: data_o = 0;
  705: data_o = 0;
  706: data_o = 0;
  707: data_o = 0;
  708: data_o = 0;
  709: data_o = 0;
  710: data_o = 1044480;
  711: data_o = 4193280;
  712: data_o = 8388352;
  713: data_o = 16777088;
  714: data_o = 33554368;
  715: data_o = 66592704;
  716: data_o = 66064352;
  717: data_o = 132122592;
  718: data_o = 132122592;
  719: data_o = 130024416;
  720: data_o = 130024432;
  721: data_o = 264242160;
  722: data_o = 264242160;
  723: data_o = 264242160;
  724: data_o = 264242160;
  725: data_o = 264242160;
  726: data_o = 2016;
  727: data_o = 2016;
  728: data_o = 2016;
  729: data_o = 4032;
  730: data_o = 4032;
  731: data_o = 8064;
  732: data_o = 16256;
  733: data_o = 16128;
  734: data_o = 32512;
  735: data_o = 65024;
  736: data_o = 130048;
  737: data_o = 260096;
  738: data_o = 258048;
  739: data_o = 516096;
  740: data_o = 1040384;
  741: data_o = 2080768;
  742: data_o = 4161536;
  743: data_o = 4128768;
  744: data_o = 8257536;
  745: data_o = 16646144;
  746: data_o = 16515072;
  747: data_o = 33030144;
  748: data_o = 66060288;
  749: data_o = 66060288;
  750: data_o = 132120576;
  751: data_o = 130023424;
  752: data_o = 264241152;
  753: data_o = 260046848;
  754: data_o = 536870904;
  755: data_o = 536870904;
  756: data_o = 536870904;
  757: data_o = 536870904;
  758: data_o = 536870904;
  759: data_o = 0;
  760: data_o = 0;
  761: data_o = 0;
  762: data_o = 0;
  763: data_o = 0;
  764: data_o = 0;
  765: data_o = 0;
  766: data_o = 0;
  767: data_o = 0;
  768: data_o = 0;
  769: data_o = 0;
  770: data_o = 0;
  771: data_o = 0;
  772: data_o = 0;
  773: data_o = 0;
  774: data_o = 2093056;
  775: data_o = 4193280;
  776: data_o = 16776704;
  777: data_o = 33554176;
  778: data_o = 33324928;
  779: data_o = 66068416;
  780: data_o = 132124608;
  781: data_o = 132122592;
  782: data_o = 130025440;
  783: data_o = 264243168;
  784: data_o = 264242144;
  785: data_o = 260047840;
  786: data_o = 260047840;
  787: data_o = 992;
  788: data_o = 992;
  789: data_o = 992;
  790: data_o = 2016;
  791: data_o = 1984;
  792: data_o = 4032;
  793: data_o = 8064;
  794: data_o = 32512;
  795: data_o = 261632;
  796: data_o = 260096;
  797: data_o = 260096;
  798: data_o = 261632;
  799: data_o = 130816;
  800: data_o = 8064;
  801: data_o = 4032;
  802: data_o = 2016;
  803: data_o = 2016;
  804: data_o = 1008;
  805: data_o = 1008;
  806: data_o = 1008;
  807: data_o = 1008;
  808: data_o = 520094704;
  809: data_o = 520094704;
  810: data_o = 528483312;
  811: data_o = 528483312;
  812: data_o = 528483312;
  813: data_o = 528483312;
  814: data_o = 264243168;
  815: data_o = 264245216;
  816: data_o = 132128704;
  817: data_o = 133726144;
  818: data_o = 67108736;
  819: data_o = 33554176;
  820: data_o = 16776704;
  821: data_o = 4192256;
  822: data_o = 507904;
  823: data_o = 0;
  824: data_o = 0;
  825: data_o = 0;
  826: data_o = 0;
  827: data_o = 0;
  828: data_o = 0;
  829: data_o = 0;
  830: data_o = 0;
  831: data_o = 0;
  832: data_o = 0;
  833: data_o = 0;
  834: data_o = 0;
  835: data_o = 0;
  836: data_o = 0;
  837: data_o = 0;
  838: data_o = 16256;
  839: data_o = 16256;
  840: data_o = 32640;
  841: data_o = 32640;
  842: data_o = 65408;
  843: data_o = 65408;
  844: data_o = 130944;
  845: data_o = 130944;
  846: data_o = 262016;
  847: data_o = 262016;
  848: data_o = 515968;
  849: data_o = 515968;
  850: data_o = 1023872;
  851: data_o = 1023872;
  852: data_o = 2039680;
  853: data_o = 2039680;
  854: data_o = 4071296;
  855: data_o = 4071296;
  856: data_o = 8134528;
  857: data_o = 8134528;
  858: data_o = 16260992;
  859: data_o = 16260992;
  860: data_o = 32513920;
  861: data_o = 32513920;
  862: data_o = 65019776;
  863: data_o = 132128640;
  864: data_o = 130031488;
  865: data_o = 264249216;
  866: data_o = 260054912;
  867: data_o = 528490368;
  868: data_o = 520101760;
  869: data_o = 1056972672;
  870: data_o = 1073741820;
  871: data_o = 1073741820;
  872: data_o = 1073741820;
  873: data_o = 1073741820;
  874: data_o = 1073741820;
  875: data_o = 8064;
  876: data_o = 8064;
  877: data_o = 8064;
  878: data_o = 8064;
  879: data_o = 8064;
  880: data_o = 8064;
  881: data_o = 8064;
  882: data_o = 8064;
  883: data_o = 8064;
  884: data_o = 8064;
  885: data_o = 8064;
  886: data_o = 8064;
  887: data_o = 0;
  888: data_o = 0;
  889: data_o = 0;
  890: data_o = 0;
  891: data_o = 0;
  892: data_o = 0;
  893: data_o = 0;
  894: data_o = 0;
  895: data_o = 0;
  896: data_o = 0;
  897: data_o = 0;
  898: data_o = 0;
  899: data_o = 0;
  900: data_o = 0;
  901: data_o = 0;
  902: data_o = 67108832;
  903: data_o = 67108832;
  904: data_o = 67108832;
  905: data_o = 67108832;
  906: data_o = 134217696;
  907: data_o = 130023424;
  908: data_o = 130023424;
  909: data_o = 130023424;
  910: data_o = 130023424;
  911: data_o = 130023424;
  912: data_o = 130023424;
  913: data_o = 130023424;
  914: data_o = 130023424;
  915: data_o = 130023424;
  916: data_o = 130023424;
  917: data_o = 130023424;
  918: data_o = 130023424;
  919: data_o = 130283520;
  920: data_o = 131071488;
  921: data_o = 132120320;
  922: data_o = 134217600;
  923: data_o = 134102976;
  924: data_o = 267915200;
  925: data_o = 266340320;
  926: data_o = 266340320;
  927: data_o = 264242144;
  928: data_o = 260047856;
  929: data_o = 1008;
  930: data_o = 1008;
  931: data_o = 1008;
  932: data_o = 1008;
  933: data_o = 1008;
  934: data_o = 1008;
  935: data_o = 1008;
  936: data_o = 1008;
  937: data_o = 528483312;
  938: data_o = 528483312;
  939: data_o = 528483312;
  940: data_o = 528484320;
  941: data_o = 528484320;
  942: data_o = 264243168;
  943: data_o = 264245184;
  944: data_o = 132128704;
  945: data_o = 133726080;
  946: data_o = 67108608;
  947: data_o = 33553920;
  948: data_o = 16776192;
  949: data_o = 8384512;
  950: data_o = 1015808;
  951: data_o = 0;
  952: data_o = 0;
  953: data_o = 0;
  954: data_o = 0;
  955: data_o = 0;
  956: data_o = 0;
  957: data_o = 0;
  958: data_o = 0;
  959: data_o = 0;
  960: data_o = 0;
  961: data_o = 0;
  962: data_o = 0;
  963: data_o = 0;
  964: data_o = 0;
  965: data_o = 0;
  966: data_o = 261120;
  967: data_o = 1048320;
  968: data_o = 2097024;
  969: data_o = 4194240;
  970: data_o = 8388544;
  971: data_o = 16650208;
  972: data_o = 16517088;
  973: data_o = 33031136;
  974: data_o = 33031152;
  975: data_o = 66061296;
  976: data_o = 66061296;
  977: data_o = 132120576;
  978: data_o = 132120576;
  979: data_o = 132120576;
  980: data_o = 130023424;
  981: data_o = 264241152;
  982: data_o = 264241152;
  983: data_o = 264370176;
  984: data_o = 264764928;
  985: data_o = 265289472;
  986: data_o = 262143872;
  987: data_o = 264241088;
  988: data_o = 268177344;
  989: data_o = 267913184;
  990: data_o = 267388896;
  991: data_o = 266339312;
  992: data_o = 266339312;
  993: data_o = 264242160;
  994: data_o = 264241648;
  995: data_o = 264241648;
  996: data_o = 264241648;
  997: data_o = 264241648;
  998: data_o = 264241648;
  999: data_o = 264241648;
  1000: data_o = 264241648;
  1001: data_o = 264241648;
  1002: data_o = 130023920;
  1003: data_o = 130024432;
  1004: data_o = 132121584;
  1005: data_o = 132121584;
  1006: data_o = 66061280;
  1007: data_o = 66062304;
  1008: data_o = 33034176;
  1009: data_o = 33431488;
  1010: data_o = 16777088;
  1011: data_o = 8388352;
  1012: data_o = 4193792;
  1013: data_o = 1047552;
  1014: data_o = 253952;
  1015: data_o = 0;
  1016: data_o = 0;
  1017: data_o = 0;
  1018: data_o = 0;
  1019: data_o = 0;
  1020: data_o = 0;
  1021: data_o = 0;
  1022: data_o = 0;
  1023: data_o = 0;
  1024: data_o = 0;
  1025: data_o = 0;
  1026: data_o = 0;
  1027: data_o = 0;
  1028: data_o = 0;
  1029: data_o = 0;
  1030: data_o = 268435440;
  1031: data_o = 268435440;
  1032: data_o = 268435440;
  1033: data_o = 268435440;
  1034: data_o = 268435440;
  1035: data_o = 1008;
  1036: data_o = 992;
  1037: data_o = 992;
  1038: data_o = 2016;
  1039: data_o = 2016;
  1040: data_o = 1984;
  1041: data_o = 1984;
  1042: data_o = 4032;
  1043: data_o = 3968;
  1044: data_o = 3968;
  1045: data_o = 3968;
  1046: data_o = 8064;
  1047: data_o = 7936;
  1048: data_o = 7936;
  1049: data_o = 16128;
  1050: data_o = 16128;
  1051: data_o = 15872;
  1052: data_o = 15872;
  1053: data_o = 32256;
  1054: data_o = 32256;
  1055: data_o = 31744;
  1056: data_o = 64512;
  1057: data_o = 64512;
  1058: data_o = 63488;
  1059: data_o = 63488;
  1060: data_o = 129024;
  1061: data_o = 129024;
  1062: data_o = 126976;
  1063: data_o = 258048;
  1064: data_o = 258048;
  1065: data_o = 258048;
  1066: data_o = 253952;
  1067: data_o = 516096;
  1068: data_o = 516096;
  1069: data_o = 507904;
  1070: data_o = 507904;
  1071: data_o = 1032192;
  1072: data_o = 1032192;
  1073: data_o = 1015808;
  1074: data_o = 2064384;
  1075: data_o = 2064384;
  1076: data_o = 2064384;
  1077: data_o = 2031616;
  1078: data_o = 4128768;
  1079: data_o = 0;
  1080: data_o = 0;
  1081: data_o = 0;
  1082: data_o = 0;
  1083: data_o = 0;
  1084: data_o = 0;
  1085: data_o = 0;
  1086: data_o = 0;
  1087: data_o = 0;
  1088: data_o = 0;
  1089: data_o = 0;
  1090: data_o = 0;
  1091: data_o = 0;
  1092: data_o = 0;
  1093: data_o = 0;
  1094: data_o = 1044480;
  1095: data_o = 4193280;
  1096: data_o = 16776704;
  1097: data_o = 33554176;
  1098: data_o = 66862976;
  1099: data_o = 66068416;
  1100: data_o = 132124608;
  1101: data_o = 130025440;
  1102: data_o = 130025440;
  1103: data_o = 264242144;
  1104: data_o = 264242144;
  1105: data_o = 264242144;
  1106: data_o = 264242144;
  1107: data_o = 264242144;
  1108: data_o = 264242144;
  1109: data_o = 264242144;
  1110: data_o = 264242144;
  1111: data_o = 130025440;
  1112: data_o = 132122560;
  1113: data_o = 65015744;
  1114: data_o = 32513920;
  1115: data_o = 33554176;
  1116: data_o = 8388096;
  1117: data_o = 2095104;
  1118: data_o = 8388096;
  1119: data_o = 33554176;
  1120: data_o = 66592640;
  1121: data_o = 132124608;
  1122: data_o = 130025440;
  1123: data_o = 264242144;
  1124: data_o = 260047856;
  1125: data_o = 528482800;
  1126: data_o = 528482808;
  1127: data_o = 528482808;
  1128: data_o = 528482808;
  1129: data_o = 528482808;
  1130: data_o = 528482808;
  1131: data_o = 528482808;
  1132: data_o = 528483312;
  1133: data_o = 528483312;
  1134: data_o = 264242160;
  1135: data_o = 266340320;
  1136: data_o = 133173216;
  1137: data_o = 133709760;
  1138: data_o = 67108736;
  1139: data_o = 33554304;
  1140: data_o = 16776704;
  1141: data_o = 4193280;
  1142: data_o = 516096;
  1143: data_o = 0;
  1144: data_o = 0;
  1145: data_o = 0;
  1146: data_o = 0;
  1147: data_o = 0;
  1148: data_o = 0;
  1149: data_o = 0;
  1150: data_o = 0;
  1151: data_o = 0;
  1152: data_o = 0;
  1153: data_o = 0;
  1154: data_o = 0;
  1155: data_o = 0;
  1156: data_o = 0;
  1157: data_o = 0;
  1158: data_o = 2088960;
  1159: data_o = 4192256;
  1160: data_o = 16776192;
  1161: data_o = 33553920;
  1162: data_o = 66879232;
  1163: data_o = 66076544;
  1164: data_o = 132128640;
  1165: data_o = 132124608;
  1166: data_o = 264243136;
  1167: data_o = 264243136;
  1168: data_o = 264243168;
  1169: data_o = 260047840;
  1170: data_o = 528483296;
  1171: data_o = 528483296;
  1172: data_o = 528483312;
  1173: data_o = 528483312;
  1174: data_o = 528483312;
  1175: data_o = 528483312;
  1176: data_o = 528483312;
  1177: data_o = 528483312;
  1178: data_o = 260047856;
  1179: data_o = 260048880;
  1180: data_o = 264243184;
  1181: data_o = 264243184;
  1182: data_o = 264245232;
  1183: data_o = 132128752;
  1184: data_o = 133185520;
  1185: data_o = 66617328;
  1186: data_o = 33553392;
  1187: data_o = 16776176;
  1188: data_o = 8381424;
  1189: data_o = 4178928;
  1190: data_o = 1008;
  1191: data_o = 992;
  1192: data_o = 2016;
  1193: data_o = 2016;
  1194: data_o = 2016;
  1195: data_o = 264245184;
  1196: data_o = 264245184;
  1197: data_o = 264245184;
  1198: data_o = 264249216;
  1199: data_o = 132136832;
  1200: data_o = 133201664;
  1201: data_o = 66649600;
  1202: data_o = 67107840;
  1203: data_o = 33553408;
  1204: data_o = 16773120;
  1205: data_o = 8380416;
  1206: data_o = 983040;
  1207: data_o = 0;
  1208: data_o = 0;
  1209: data_o = 0;
  1210: data_o = 0;
  1211: data_o = 0;
  1212: data_o = 0;
  1213: data_o = 0;
  1214: data_o = 0;
  1215: data_o = 0;
  default: data_o = 'X;
endcase
endmodule
