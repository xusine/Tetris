module memory_str_next#(
  parameter integer width_p
  parameter integer depth_p
)(
  input [depth_p-1:0] addr_i
  ,output logic [width_p-1:0] data_o
);
always unique case(addr_i)
  0: data_o = 0;
  1: data_o = 0;
  2: data_o = 0;
  3: data_o = 0;
  4: data_o = 0;
  5: data_o = 0;
  6: data_o = 0;
  7: data_o = 0;
  8: data_o = 0;
  9: data_o = 0;
  10: data_o = 0;
  11: data_o = 2143290367;
  12: data_o = 2145387519;
  13: data_o = 132120636;
  14: data_o = 133169208;
  15: data_o = 133169208;
  16: data_o = 133693496;
  17: data_o = 133693496;
  18: data_o = 133955640;
  19: data_o = 134086712;
  20: data_o = 134086712;
  21: data_o = 134152248;
  22: data_o = 125763640;
  23: data_o = 125796408;
  24: data_o = 121602104;
  25: data_o = 121618488;
  26: data_o = 119521336;
  27: data_o = 118480952;
  28: data_o = 118480952;
  29: data_o = 117960760;
  30: data_o = 117960760;
  31: data_o = 117700664;
  32: data_o = 117700664;
  33: data_o = 117570616;
  34: data_o = 117570616;
  35: data_o = 117505592;
  36: data_o = 117505592;
  37: data_o = 117473080;
  38: data_o = 117473208;
  39: data_o = 117456824;
  40: data_o = 117456888;
  41: data_o = 117448696;
  42: data_o = 117448696;
  43: data_o = 117444600;
  44: data_o = 117444600;
  45: data_o = 117442552;
  46: data_o = 117441528;
  47: data_o = 117441528;
  48: data_o = 117441016;
  49: data_o = 117441016;
  50: data_o = 117440760;
  51: data_o = 117440760;
  52: data_o = 125829240;
  53: data_o = 2146435192;
  54: data_o = 2146435128;
  55: data_o = 0;
  56: data_o = 0;
  57: data_o = 0;
  58: data_o = 0;
  59: data_o = 0;
  60: data_o = 0;
  61: data_o = 0;
  62: data_o = 0;
  63: data_o = 0;
  64: data_o = 0;
  65: data_o = 0;
  66: data_o = 0;
  67: data_o = 0;
  68: data_o = 0;
  69: data_o = 0;
  70: data_o = 0;
  71: data_o = 0;
  72: data_o = 0;
  73: data_o = 0;
  74: data_o = 0;
  75: data_o = 0;
  76: data_o = 0;
  77: data_o = 0;
  78: data_o = 0;
  79: data_o = 0;
  80: data_o = 0;
  81: data_o = 0;
  82: data_o = 0;
  83: data_o = 0;
  84: data_o = 0;
  85: data_o = 0;
  86: data_o = 0;
  87: data_o = 0;
  88: data_o = 0;
  89: data_o = 523264;
  90: data_o = 2096896;
  91: data_o = 8388544;
  92: data_o = 16719840;
  93: data_o = 33294320;
  94: data_o = 33031152;
  95: data_o = 66060792;
  96: data_o = 132121080;
  97: data_o = 132121080;
  98: data_o = 132120828;
  99: data_o = 264241404;
  100: data_o = 264241404;
  101: data_o = 264241404;
  102: data_o = 268435452;
  103: data_o = 268435452;
  104: data_o = 268435452;
  105: data_o = 264241152;
  106: data_o = 264241152;
  107: data_o = 264241152;
  108: data_o = 264241152;
  109: data_o = 132120576;
  110: data_o = 132120696;
  111: data_o = 132120696;
  112: data_o = 66060536;
  113: data_o = 66585072;
  114: data_o = 33293280;
  115: data_o = 16715744;
  116: data_o = 8388544;
  117: data_o = 4194048;
  118: data_o = 523264;
  119: data_o = 0;
  120: data_o = 0;
  121: data_o = 0;
  122: data_o = 0;
  123: data_o = 0;
  124: data_o = 0;
  125: data_o = 0;
  126: data_o = 0;
  127: data_o = 0;
  128: data_o = 0;
  129: data_o = 0;
  130: data_o = 0;
  131: data_o = 0;
  132: data_o = 0;
  133: data_o = 0;
  134: data_o = 0;
  135: data_o = 0;
  136: data_o = 0;
  137: data_o = 0;
  138: data_o = 0;
  139: data_o = 0;
  140: data_o = 0;
  141: data_o = 0;
  142: data_o = 0;
  143: data_o = 0;
  144: data_o = 0;
  145: data_o = 0;
  146: data_o = 0;
  147: data_o = 0;
  148: data_o = 0;
  149: data_o = 0;
  150: data_o = 0;
  151: data_o = 0;
  152: data_o = 0;
  153: data_o = 268386300;
  154: data_o = 268386300;
  155: data_o = 33294304;
  156: data_o = 16517056;
  157: data_o = 16648064;
  158: data_o = 8261504;
  159: data_o = 8331008;
  160: data_o = 4169216;
  161: data_o = 2080256;
  162: data_o = 2096128;
  163: data_o = 1047552;
  164: data_o = 1046528;
  165: data_o = 520192;
  166: data_o = 520192;
  167: data_o = 258048;
  168: data_o = 260096;
  169: data_o = 523264;
  170: data_o = 1047552;
  171: data_o = 1048064;
  172: data_o = 2063872;
  173: data_o = 4095744;
  174: data_o = 4079360;
  175: data_o = 8134528;
  176: data_o = 7872384;
  177: data_o = 16256960;
  178: data_o = 32509920;
  179: data_o = 32507872;
  180: data_o = 133171192;
  181: data_o = 1073496062;
  182: data_o = 1073496062;
  183: data_o = 0;
  184: data_o = 0;
  185: data_o = 0;
  186: data_o = 0;
  187: data_o = 0;
  188: data_o = 0;
  189: data_o = 0;
  190: data_o = 0;
  191: data_o = 0;
  192: data_o = 0;
  193: data_o = 0;
  194: data_o = 0;
  195: data_o = 0;
  196: data_o = 0;
  197: data_o = 0;
  198: data_o = 0;
  199: data_o = 0;
  200: data_o = 0;
  201: data_o = 0;
  202: data_o = 0;
  203: data_o = 0;
  204: data_o = 0;
  205: data_o = 0;
  206: data_o = 0;
  207: data_o = 491520;
  208: data_o = 491520;
  209: data_o = 491520;
  210: data_o = 491520;
  211: data_o = 1015808;
  212: data_o = 1015808;
  213: data_o = 1015808;
  214: data_o = 2064384;
  215: data_o = 4161536;
  216: data_o = 16744448;
  217: data_o = 268435424;
  218: data_o = 268435424;
  219: data_o = 268435424;
  220: data_o = 2064384;
  221: data_o = 2064384;
  222: data_o = 2064384;
  223: data_o = 2064384;
  224: data_o = 2064384;
  225: data_o = 2064384;
  226: data_o = 2064384;
  227: data_o = 2064384;
  228: data_o = 2064384;
  229: data_o = 2064384;
  230: data_o = 2064384;
  231: data_o = 2064384;
  232: data_o = 2064384;
  233: data_o = 2064384;
  234: data_o = 2064384;
  235: data_o = 2064384;
  236: data_o = 2064384;
  237: data_o = 2064384;
  238: data_o = 2064440;
  239: data_o = 2064504;
  240: data_o = 2064504;
  241: data_o = 2081008;
  242: data_o = 1032432;
  243: data_o = 1041376;
  244: data_o = 524256;
  245: data_o = 262080;
  246: data_o = 130816;
  247: data_o = 0;
  248: data_o = 0;
  249: data_o = 0;
  250: data_o = 0;
  251: data_o = 0;
  252: data_o = 0;
  253: data_o = 0;
  254: data_o = 0;
  255: data_o = 0;
  default: data_o = 'X;
endcase
endmodule
