package tetris;

typedef enum {eNOP, eStart, eNewTile, eRotate, eDown, eLeft, eRight} tile_opcode_e;

endpackage