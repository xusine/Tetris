package layout_parameters;

typedef struct {
  integer x_m
  ,integer y_m
} ppoint_t;

parameter ppoint_t str_score_p;

parameter ppoint_t score_pos_p;

parameter ppoint_t str_next_p;

parameter ppoint_t next_block_p;
parameter ppoint_t next_block_size_p;

parameter ppoint_t game_board_p;


endpackage

